module rv32i(
    //Entradas
    // - No estoy seguro, creo que de la memoria

    //Salidas
    // - Same
);


endmodule